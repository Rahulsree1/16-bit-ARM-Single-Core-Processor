module Imem(adr,rst,Imaout);
    input [4:0] adr;
    input [0:0] rst;
    
    output [15:0] Imaout;

    reg [15:0] mem [32:0];


    assign Imaout = (rst == 1'b0) ? 16'b0000000000000000 : mem[adr];

    initial begin

        // LDR
        mem[0] = {{5'b00000},{3'b111},{3'b001},{3'b000},{2'b01}};
        //mem[1] = {{5'b00001},{3'b111},{3'b010},{3'b000},{2'b01}};


        // R-type Instructions ADD SUB AND OR NOT XOR
        // mem[2] = {{2'b00},{3'b010},{3'b001},{3'b011},{3'b000},{2'b00}};
        // mem[3] = {{2'b00},{3'b010},{3'b001},{3'b100},{3'b001},{2'b00}};
        // mem[4] = {{2'b00},{3'b001},{3'b011},{3'b010},{3'b010},{2'b00}};
        // mem[5] = {{2'b00},{3'b001},{3'b011},{3'b010},{3'b011},{2'b00}};
        // mem[6] = {{2'b00},{3'b001},{3'b011},{3'b010},{3'b100},{2'b00}};
        // mem[7] = {{2'b00},{3'b001},{3'b011},{3'b010},{3'b101},{2'b00}};


        

        // I - type LOAD 
        // STORE
        // mem[8] = {{5'b00000},{3'b111},{3'b110},{3'b000},{2'b11}};   // address src
        // mem[1] = {{5'b00000},{3'b010},{3'b111},{3'b000},{2'b01}};


        // B - type
        //mem[0] = {{5'b00010},{3'b010},{3'b001},{3'b000},{2'b10}};

        // mem[5'b00010] = {{2'b00},{3'b001},{3'b110},{3'b010},{3'b000},{2'b00}};

        //Function Call

        // mem[0] = {{2'b00},{3'b001},{3'b011},{3'b110},{3'b000},{2'b00}};
        // mem[1] = {{6'b000000},{5'b01010},{3'b110},{2'b11}};// function call
        // mem[2] = {{2'b00},{3'b001},{3'b011},{3'b110},{3'b000},{2'b00}}; 
        
        
        //function
        // mem[5'b01010] = {{5'b00000},{3'b010},{3'b111},{3'b000},{2'b01}};
        // mem[5'b01011] = {{6'b111111},{5'b01010},{3'b111},{2'b11}}; //function call return

        // mem[0] = {{2'b00},{3'b001},{3'b011},{3'b110},{3'b000},{2'b00}};
        // mem[1] = {{2'b00},{3'b001},{3'b011},{3'b110},{3'b000},{2'b00}};
        // mem[2] = {16{1'b1}};
        
    end


endmodule






 
